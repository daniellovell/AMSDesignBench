Vin vin 0 AC 1

Rin vin nsum ?
Rfb1 z nsum ?
Rfb2 y nsum ?
XU1 u nsum 0 OPAMP

Rint1 u n2 ?
Cint1 y n2 ?
XU2 y n2 0 OPAMP

Rint2 y n3 ?
Cint2 z n3 ?
XU3 z n3 0 OPAMP

Rload y 0 ?

.end
