Vin vin 0 AC 1
L1 vin vout BLANK
R1 vout 0 BLANK
Rload vout 0 BLANK

.end
