* Working SKY130 Gm/ID Test using .print
.option scale=1.0u

* Define required slope parameters
.param sky130_fd_pr__nfet_01v8__toxe_slope = 0
.param sky130_fd_pr__nfet_01v8__vth0_slope = 0  
.param sky130_fd_pr__nfet_01v8__vth0_slope1 = 0
.param sky130_fd_pr__nfet_01v8__voff_slope = 0
.param sky130_fd_pr__nfet_01v8__nfactor_slope = 0
.param sky130_fd_pr__nfet_01v8__lint_diff = 0
.param sky130_fd_pr__nfet_01v8__wint_diff = 0

* Include SKY130 NFET model
.include cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice

* Test circuit
Vdd vdd 0 DC 1.8
Vss vss 0 DC 0
Vgs vgs 0 DC 0.6

* NFET: Drain=vdd, Gate=vgs, Source=vss, Bulk=vss
XM1 vdd vgs vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1

* DC sweep
.dc Vgs 0 1.2 0.05

* Print device parameters
.print dc v(vgs) @xm1.msky130_fd_pr__nfet_01v8[id] @xm1.msky130_fd_pr__nfet_01v8[gm] @xm1.msky130_fd_pr__nfet_01v8[gds]

.end

