Vin vin 0 AC 1
C1 vin n1 BLANK
R2 vout n1 BLANK
C2 vout n1 BLANK
R3 n1 0 BLANK
XU1 vout n1 0 OPAMP
Rload vout 0 BLANK

.end
