Vin vin 0 AC 1
R1 vin nA BLANK
R2 nA vout BLANK
Cmid nA 0 BLANK
C1 vin nB BLANK
C2 nB vout BLANK
Rmid nB 0 BLANK
Rload vout 0 BLANK

.end
