Vin vin 0 AC 1
C1 vin n1 BLANK
C2 n1 vout BLANK
R1 n1 0 BLANK
R2 vout 0 BLANK
XU1 vout vout n1 OPAMP
Rload vout 0 BLANK

.end
