Vin vin 0 AC 1
R1A vin n1 BLANK
R2A n1 v1 BLANK
C1A n1 0 BLANK
C2A v1 n1 BLANK
XU1 v1 n1i v1 OPAMP
RG1 n1i 0 BLANK
RF1 v1 n1i BLANK

 
R1B v1 n2 BLANK
R2B n2 vout BLANK
C1B n2 0 BLANK
C2B vout n2 BLANK
XU2 vout n2i vout OPAMP
RG2 n2i 0 BLANK
RF2 vout n2i BLANK

Rload vout 0 BLANK

.end
