Vin vin 0 AC 1

Rin vin nsum ?
Rfb1 z nsum ?
Rfb2 vout nsum ?
XU1 u nsum 0 OPAMP

Rint1 u n2 ?
Cint1 vout n2 ?
XU2 vout n2 0 OPAMP

Rint2 vout n3 ?
Cint2 z n3 ?
XU3 z n3 0 OPAMP

Rload vout 0 ?

.end
