Vin vin 0 AC 1
R1 vin npos BLANK
C1 npos 0 BLANK
R2 vin nneg BLANK
R3 vout nneg BLANK
XU1 vout nneg npos OPAMP
Rload vout 0 BLANK

.end
