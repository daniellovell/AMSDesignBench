Vin vin 0 AC 1
R1A vin n1 ?
R2A n1 v1 ?
C1A n1 0 ?
C2A v1 n1 ?
XU1 v1 n1i v1 OPAMP
RG1 n1i 0 ?
RF1 v1 n1i ?

 
R1B v1 n2 ?
R2B n2 vout ?
C1B n2 0 ?
C2B vout n2 ?
XU2 vout n2i vout OPAMP
RG2 n2i 0 ?
RF2 vout n2i ?

Rload vout 0 ?

.end
