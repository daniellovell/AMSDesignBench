Vin vin 0 AC 1
L1 vin vout ?
R1 vout 0 ?
Rload vout 0 ?

.end
