Vin vin 0 AC 1
R1 vin npos ?
C1 npos 0 ?
R2 vin nneg ?
R3 vout nneg ?
XU1 vout nneg npos OPAMP
Rload vout 0 ?

.end
