Vin vin 0 AC 1
R1 vin n1 ?
C1 n1 nneg ?
C2 vout n2 ?
R2 n2 nneg ?
XU1 vout nneg 0 OPAMP
Rload vout 0 ?

.end
