Vin vin 0 AC 1
C1 vin n1 ?
R2 vout n1 ?
C2 vout n1 ?
R3 n1 0 ?
XU1 vout n1 0 OPAMP
Rload vout 0 ?

.end
