Vin vin 0 AC 1

Rin vin nsum BLANK
Rfb1 z nsum BLANK
Rfb2 vout nsum BLANK
XU1 u nsum 0 OPAMP

Rint1 u n2 BLANK
Cint1 vout n2 BLANK
XU2 vout n2 0 OPAMP

Rint2 vout n3 BLANK
Cint2 z n3 BLANK
XU3 z n3 0 OPAMP

Rload vout 0 BLANK

.end
