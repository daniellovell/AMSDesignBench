Vin vin 0 AC 1
R1 vin nA ?
R2 nA vout ?
Cmid nA 0 ?
C1 vin nB ?
C2 nB vout ?
Rmid nB 0 ?
Rload vout 0 ?

.end
