Vin vin 0 AC 1
C1 vin n1 ?
C2 n1 vout ?
R1 n1 0 ?
R2 vout 0 ?
XU1 vout vout n1 OPAMP
Rload vout 0 ?

.end
