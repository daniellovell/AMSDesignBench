* Noninverting Voltage Amplifier with Resistive Feedback
subckt opamp in_n in_p out
	* opamp implementation
ends opamp
XU1 N001 S_in S_out opamp Aol=100K GBW=10Meg
R1 0 N001 R
R2 S_out N001 R
.backanno
.end

